package axis_fifo_pkg_prm;

    parameter AXI_DATA_WIDTH = 32;
    parameter AXI_DATA_DEPTH = 1024;

endpackage