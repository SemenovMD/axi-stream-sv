package axis_uart_pkg_prm;

    parameter AXI_DATA_WIDTH    = 32;

    parameter CLOCK             = 100_000_000;

    parameter BAUD_RATE         = 115_200;
    parameter DATA_BITS         = 8;
    parameter STOP_BITS         = 1;
    parameter PARITY_BITS       = 0;

endpackage