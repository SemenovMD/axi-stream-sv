package axis_crc32_mpeg2_pkg_prm;

    parameter AXI_DATA_WIDTH = 32;
    parameter INIT_CRC       = 32'hFFFF_FFFF;
    parameter POLY_CRC       = 32'h04C1_1DB7;

endpackage
