package pkg_tb;

    parameter AXI_DATA_WIDTH = 32;
    parameter AXI_DATA_DEPTH = 32;

    parameter AXI_TRAN_MIN_DELAY = 2;
    parameter AXI_TRAN_MAX_DELAY = 17;

    parameter AXI_TRAN_MAX_WAIT = 150;

endpackage