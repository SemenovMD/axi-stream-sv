package axis_converter_lite_pkg_prm;

    parameter AXI_DATA_WIDTH    = 32;
    parameter AXI_ADDR_WIDTH    = 32;

    parameter AXI_ADDR          = 32'h0000_0001;

endpackage