package axis_uart_pkg_tb;

    import axis_uart_pkg_prm::*;

    parameter AXI_TRAN_MIN_DELAY = 2;
    parameter AXI_TRAN_MAX_DELAY = 17;

    parameter UART_RX_MIN_DELAY = 5;
    parameter UART_RX_MAX_DELAY = 20;

endpackage